module TopLevel();


endmodule: TopLevel