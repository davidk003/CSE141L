module MemoryController(
    input logic regToReg,
    input logic regToMem,
    input logic memToReg,
    input logic [7:0] regData,
    input logic [7:0] ALUdata,
    input logic [7:0] address
    output logic 
);

always_comb begin
    if (regToReg) begin
       
    end
    else if (regToMem) begin
        
    end
end



endmodule