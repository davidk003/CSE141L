module ALUout(
    input  writeBack,
    input logic [7:0] Rslt,
    input logic [2:0] reg
    input logic [7:0] dataOut
);

endmodule