module ALUInMux ( 
	input logic writeBack,
	input logic [1:0] reg1,
	input logic [1:0] reg2,
	input logic [2:0] Aluop,
	output logic [7:0] op1,
	output logic [7:0] op2
   );
   //Mux input for ALU

always_comb begin
	
end
endmodule
